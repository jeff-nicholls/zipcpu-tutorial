//////////////////////////////////////////////////////////////////////////////////
// thruwire.sv
// Jeff Nicholls
// 2024
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps
`default_nettype none

module thruwire(
    input wire SW,
    output wire LED
    );
    
    assign LED = SW;
        
endmodule
